module discordv