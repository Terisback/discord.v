module structs

pub struct Member {
	
}