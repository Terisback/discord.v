module types

// Intent type for gateway connection
pub type Intent = u16

// Permission type
pub type Permission = int