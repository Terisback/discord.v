module discordv

// Constants for general managment
pub const (
	create_instant_invite = Permission(0x00000001)
	kick_members          = Permission(0x00000002)
	ban_members           = Permission(0x00000004)
	administrator         = Permission(0x00000008)
	manage_channels       = Permission(0x00000010)
	manage_guild          = Permission(0x00000020)
	add_reactions         = Permission(0x00000040)
	view_audit_log        = Permission(0x00000080)
	priority_speaker      = Permission(0x00000100)
	stream                = Permission(0x00000200)
	view_channel          = Permission(0x00000400)
	send_messages         = Permission(0x00000800)
	send_tts_messages     = Permission(0x00001000)
	manage_messages       = Permission(0x00002000)
	embed_links           = Permission(0x00004000)
	attach_files          = Permission(0x00008000)
	read_message_history  = Permission(0x00010000)
	mention_everyone      = Permission(0x00020000)
	use_external_emojis   = Permission(0x00040000)
	view_guild_insights   = Permission(0x00080000)
	connect               = Permission(0x00100000)
	speak                 = Permission(0x00200000)
	mute_members          = Permission(0x00400000)
	deafen_members        = Permission(0x00800000)
	move_members          = Permission(0x01000000)
	use_vad               = Permission(0x02000000)
	change_nickname       = Permission(0x04000000)
	manage_nicknames      = Permission(0x08000000)
	manage_roles          = Permission(0x10000000)
	manage_webhooks       = Permission(0x20000000)
	manage_emojis         = Permission(0x40000000)
)
