module structs

pub struct Resumed {} // lul, it's empty