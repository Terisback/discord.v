module structs

pub struct Channel {
	
}