module types

pub type Permission = int