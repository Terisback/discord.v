module packets

// Websocket Hello packet data
pub struct Hello {
pub:
	heartbeat_interval u64
}
