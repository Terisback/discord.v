module rest

struct RateLimit {
	// TODO
}