module structs

pub struct Attachment {
	
}