module structs

pub struct User {
	
}