module structs

pub struct Reconnect {
pub:
	resumed bool
}