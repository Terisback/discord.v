module structs

pub struct Reaction {
	count int
	me bool
	emoji Emoji
}