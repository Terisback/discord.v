module discordv

import discordv.types

// Constants for the different bit offsets of intents
pub const (
	guilds                   = types.Intent(1 << 0)
	guild_members            = types.Intent(1 << 1)
	guild_bans               = types.Intent(1 << 2)
	guild_emojis             = types.Intent(1 << 3)
	guild_integrations       = types.Intent(1 << 4)
	guild_webhooks           = types.Intent(1 << 5)
	guild_invites            = types.Intent(1 << 6)
	guild_voice_states       = types.Intent(1 << 7)
	guild_precenses          = types.Intent(1 << 8)
	guild_messages           = types.Intent(1 << 9)
	guild_message_reactions  = types.Intent(1 << 10)
	guild_message_typing     = types.Intent(1 << 11)
	direct_messages          = types.Intent(1 << 12)
	direct_message_reactions = types.Intent(1 << 13)
	direct_message_typing    = types.Intent(1 << 14)
	all_allowed              = types.Intent(32509)
	all                      = types.Intent(32767)
)

// Constants for general managment
pub const (
	create_instant_invite = types.Permission(0x00000001)
	kick_members          = types.Permission(0x00000002)
	ban_members           = types.Permission(0x00000004)
	administrator         = types.Permission(0x00000008)
	manage_channels       = types.Permission(0x00000010)
	manage_guild          = types.Permission(0x00000020)
	add_reactions         = types.Permission(0x00000040)
	view_audit_log        = types.Permission(0x00000080)
	priority_speaker      = types.Permission(0x00000100)
	stream                = types.Permission(0x00000200)
	view_channel          = types.Permission(0x00000400)
	send_messages         = types.Permission(0x00000800)
	send_tts_messages     = types.Permission(0x00001000)
	manage_messages       = types.Permission(0x00002000)
	embed_links           = types.Permission(0x00004000)
	attach_files          = types.Permission(0x00008000)
	read_message_history  = types.Permission(0x00010000)
	mention_everyone      = types.Permission(0x00020000)
	use_external_emojis   = types.Permission(0x00040000)
	view_guild_insights   = types.Permission(0x00080000)
	connect               = types.Permission(0x00100000)
	speak                 = types.Permission(0x00200000)
	mute_members          = types.Permission(0x00400000)
	deafen_members        = types.Permission(0x00800000)
	move_members          = types.Permission(0x01000000)
	use_vad               = types.Permission(0x02000000)
	change_nickname       = types.Permission(0x04000000)
	manage_nicknames      = types.Permission(0x08000000)
	manage_roles          = types.Permission(0x10000000)
	manage_webhooks       = types.Permission(0x20000000)
	manage_emojis         = types.Permission(0x40000000)
)
