module structs

pub struct File {
pub mut:
	filename string
	data []byte
}