module structs

pub struct Reaction {
	
}