module client

struct RateLimit {
	
}