module structs

pub struct Embed {
	
}