module types

pub type Intent = u16